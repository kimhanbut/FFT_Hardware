`timescale 1ns / 1ps

module cos_rom (
    input  logic        clk,
    input  logic [8:0]  addr,              // 9-bit address (0 ~ 496, 16단위)
    output logic [8:0]  data [0:15]        // 16개의 9-bit 병렬 출력
);

  logic [8:0] mem [0:511];

  // 합성 가능한 방식: 직접 초기화
  // *** 주의: 아래는 예시이며, 실제로는 512개의 데이터가 모두 필요합니다 ***
  initial begin
    mem[0]  = 9'b000111111;
    mem[1]  = 9'b001000000;
    mem[2]  = 9'b001000000;
    mem[3]  = 9'b001000000;
    mem[4]  = 9'b001000000;
    mem[5]  = 9'b001000000;
    mem[6]  = 9'b001000000;
    mem[7]  = 9'b001000000;
    mem[8]  = 9'b001000000;
    mem[9]  = 9'b001000000;
    mem[10]  = 9'b001000000;
    mem[11]  = 9'b000111111;
    mem[12]  = 9'b000111111;
    mem[13]  = 9'b000111111;
    mem[14]  = 9'b000111111;
    mem[15]  = 9'b000111111;
    mem[16]  = 9'b000111111;
    mem[17]  = 9'b000111111;
    mem[18]  = 9'b000111110;
    mem[19]  = 9'b000111110;
    mem[20]  = 9'b000111110;
    mem[21]  = 9'b000111110;
    mem[22]  = 9'b000111110;
    mem[23]  = 9'b000111101;
    mem[24]  = 9'b000111101;
    mem[25]  = 9'b000111101;
    mem[26]  = 9'b000111101;
    mem[27]  = 9'b000111101;
    mem[28]  = 9'b000111100;
    mem[29]  = 9'b000111100;
    mem[30]  = 9'b000111100;
    mem[31]  = 9'b000111011;
    mem[32]  = 9'b000111011;
    mem[33]  = 9'b000111011;
    mem[34]  = 9'b000111011;
    mem[35]  = 9'b000111010;
    mem[36]  = 9'b000111010;
    mem[37]  = 9'b000111010;
    mem[38]  = 9'b000111001;
    mem[39]  = 9'b000111001;
    mem[40]  = 9'b000111000;
    mem[41]  = 9'b000111000;
    mem[42]  = 9'b000111000;
    mem[43]  = 9'b000110111;
    mem[44]  = 9'b000110111;
    mem[45]  = 9'b000110110;
    mem[46]  = 9'b000110110;
    mem[47]  = 9'b000110110;
    mem[48]  = 9'b000110101;
    mem[49]  = 9'b000110101;
    mem[50]  = 9'b000110100;
    mem[51]  = 9'b000110100;
    mem[52]  = 9'b000110011;
    mem[53]  = 9'b000110011;
    mem[54]  = 9'b000110010;
    mem[55]  = 9'b000110010;
    mem[56]  = 9'b000110001;
    mem[57]  = 9'b000110001;
    mem[58]  = 9'b000110000;
    mem[59]  = 9'b000110000;
    mem[60]  = 9'b000101111;
    mem[61]  = 9'b000101111;
    mem[62]  = 9'b000101110;
    mem[63]  = 9'b000101110;
    mem[64]  = 9'b000101101;
    mem[65]  = 9'b000101101;
    mem[66]  = 9'b000101100;
    mem[67]  = 9'b000101100;
    mem[68]  = 9'b000101011;
    mem[69]  = 9'b000101010;
    mem[70]  = 9'b000101010;
    mem[71]  = 9'b000101001;
    mem[72]  = 9'b000101001;
    mem[73]  = 9'b000101000;
    mem[74]  = 9'b000100111;
    mem[75]  = 9'b000100111;
    mem[76]  = 9'b000100110;
    mem[77]  = 9'b000100101;
    mem[78]  = 9'b000100101;
    mem[79]  = 9'b000100100;
    mem[80]  = 9'b000100100;
    mem[81]  = 9'b000100011;
    mem[82]  = 9'b000100010;
    mem[83]  = 9'b000100010;
    mem[84]  = 9'b000100001;
    mem[85]  = 9'b000100000;
    mem[86]  = 9'b000100000;
    mem[87]  = 9'b000011111;
    mem[88]  = 9'b000011110;
    mem[89]  = 9'b000011101;
    mem[90]  = 9'b000011101;
    mem[91]  = 9'b000011100;
    mem[92]  = 9'b000011011;
    mem[93]  = 9'b000011011;
    mem[94]  = 9'b000011010;
    mem[95]  = 9'b000011001;
    mem[96]  = 9'b000011000;
    mem[97]  = 9'b000011000;
    mem[98]  = 9'b000010111;
    mem[99]  = 9'b000010110;
    mem[100]  = 9'b000010110;
    mem[101]  = 9'b000010101;
    mem[102]  = 9'b000010100;
    mem[103]  = 9'b000010011;
    mem[104]  = 9'b000010011;
    mem[105]  = 9'b000010010;
    mem[106]  = 9'b000010001;
    mem[107]  = 9'b000010000;
    mem[108]  = 9'b000010000;
    mem[109]  = 9'b000001111;
    mem[110]  = 9'b000001110;
    mem[111]  = 9'b000001101;
    mem[112]  = 9'b000001100;
    mem[113]  = 9'b000001100;
    mem[114]  = 9'b000001011;
    mem[115]  = 9'b000001010;
    mem[116]  = 9'b000001001;
    mem[117]  = 9'b000001001;
    mem[118]  = 9'b000001000;
    mem[119]  = 9'b000000111;
    mem[120]  = 9'b000000110;
    mem[121]  = 9'b000000101;
    mem[122]  = 9'b000000101;
    mem[123]  = 9'b000000100;
    mem[124]  = 9'b000000011;
    mem[125]  = 9'b000000010;
    mem[126]  = 9'b000000010;
    mem[127]  = 9'b000000001;
    mem[128]  = 9'b000000000;
    mem[129]  = 9'b111111111;
    mem[130]  = 9'b111111110;
    mem[131]  = 9'b111111110;
    mem[132]  = 9'b111111101;
    mem[133]  = 9'b111111100;
    mem[134]  = 9'b111111011;
    mem[135]  = 9'b111111011;
    mem[136]  = 9'b111111010;
    mem[137]  = 9'b111111001;
    mem[138]  = 9'b111111000;
    mem[139]  = 9'b111110111;
    mem[140]  = 9'b111110111;
    mem[141]  = 9'b111110110;
    mem[142]  = 9'b111110101;
    mem[143]  = 9'b111110100;
    mem[144]  = 9'b111110100;
    mem[145]  = 9'b111110011;
    mem[146]  = 9'b111110010;
    mem[147]  = 9'b111110001;
    mem[148]  = 9'b111110000;
    mem[149]  = 9'b111110000;
    mem[150]  = 9'b111101111;
    mem[151]  = 9'b111101110;
    mem[152]  = 9'b111101101;
    mem[153]  = 9'b111101101;
    mem[154]  = 9'b111101100;
    mem[155]  = 9'b111101011;
    mem[156]  = 9'b111101010;
    mem[157]  = 9'b111101010;
    mem[158]  = 9'b111101001;
    mem[159]  = 9'b111101000;
    mem[160]  = 9'b111101000;
    mem[161]  = 9'b111100111;
    mem[162]  = 9'b111100110;
    mem[163]  = 9'b111100101;
    mem[164]  = 9'b111100101;
    mem[165]  = 9'b111100100;
    mem[166]  = 9'b111100011;
    mem[167]  = 9'b111100011;
    mem[168]  = 9'b111100010;
    mem[169]  = 9'b111100001;
    mem[170]  = 9'b111100000;
    mem[171]  = 9'b111100000;
    mem[172]  = 9'b111011111;
    mem[173]  = 9'b111011110;
    mem[174]  = 9'b111011110;
    mem[175]  = 9'b111011101;
    mem[176]  = 9'b111011100;
    mem[177]  = 9'b111011100;
    mem[178]  = 9'b111011011;
    mem[179]  = 9'b111011011;
    mem[180]  = 9'b111011010;
    mem[181]  = 9'b111011001;
    mem[182]  = 9'b111011001;
    mem[183]  = 9'b111011000;
    mem[184]  = 9'b111010111;
    mem[185]  = 9'b111010111;
    mem[186]  = 9'b111010110;
    mem[187]  = 9'b111010110;
    mem[188]  = 9'b111010101;
    mem[189]  = 9'b111010100;
    mem[190]  = 9'b111010100;
    mem[191]  = 9'b111010011;
    mem[192]  = 9'b111010011;
    mem[193]  = 9'b111010010;
    mem[194]  = 9'b111010010;
    mem[195]  = 9'b111010001;
    mem[196]  = 9'b111010001;
    mem[197]  = 9'b111010000;
    mem[198]  = 9'b111010000;
    mem[199]  = 9'b111001111;
    mem[200]  = 9'b111001111;
    mem[201]  = 9'b111001110;
    mem[202]  = 9'b111001110;
    mem[203]  = 9'b111001101;
    mem[204]  = 9'b111001101;
    mem[205]  = 9'b111001100;
    mem[206]  = 9'b111001100;
    mem[207]  = 9'b111001011;
    mem[208]  = 9'b111001011;
    mem[209]  = 9'b111001010;
    mem[210]  = 9'b111001010;
    mem[211]  = 9'b111001010;
    mem[212]  = 9'b111001001;
    mem[213]  = 9'b111001001;
    mem[214]  = 9'b111001000;
    mem[215]  = 9'b111001000;
    mem[216]  = 9'b111001000;
    mem[217]  = 9'b111000111;
    mem[218]  = 9'b111000111;
    mem[219]  = 9'b111000110;
    mem[220]  = 9'b111000110;
    mem[221]  = 9'b111000110;
    mem[222]  = 9'b111000101;
    mem[223]  = 9'b111000101;
    mem[224]  = 9'b111000101;
    mem[225]  = 9'b111000101;
    mem[226]  = 9'b111000100;
    mem[227]  = 9'b111000100;
    mem[228]  = 9'b111000100;
    mem[229]  = 9'b111000011;
    mem[230]  = 9'b111000011;
    mem[231]  = 9'b111000011;
    mem[232]  = 9'b111000011;
    mem[233]  = 9'b111000011;
    mem[234]  = 9'b111000010;
    mem[235]  = 9'b111000010;
    mem[236]  = 9'b111000010;
    mem[237]  = 9'b111000010;
    mem[238]  = 9'b111000010;
    mem[239]  = 9'b111000001;
    mem[240]  = 9'b111000001;
    mem[241]  = 9'b111000001;
    mem[242]  = 9'b111000001;
    mem[243]  = 9'b111000001;
    mem[244]  = 9'b111000001;
    mem[245]  = 9'b111000001;
    mem[246]  = 9'b111000000;
    mem[247]  = 9'b111000000;
    mem[248]  = 9'b111000000;
    mem[249]  = 9'b111000000;
    mem[250]  = 9'b111000000;
    mem[251]  = 9'b111000000;
    mem[252]  = 9'b111000000;
    mem[253]  = 9'b111000000;
    mem[254]  = 9'b111000000;
    mem[255]  = 9'b111000000;
    mem[256]  = 9'b111000000;
    mem[257]  = 9'b111000000;
    mem[258]  = 9'b111000000;
    mem[259]  = 9'b111000000;
    mem[260]  = 9'b111000000;
    mem[261]  = 9'b111000000;
    mem[262]  = 9'b111000000;
    mem[263]  = 9'b111000000;
    mem[264]  = 9'b111000000;
    mem[265]  = 9'b111000000;
    mem[266]  = 9'b111000000;
    mem[267]  = 9'b111000001;
    mem[268]  = 9'b111000001;
    mem[269]  = 9'b111000001;
    mem[270]  = 9'b111000001;
    mem[271]  = 9'b111000001;
    mem[272]  = 9'b111000001;
    mem[273]  = 9'b111000001;
    mem[274]  = 9'b111000010;
    mem[275]  = 9'b111000010;
    mem[276]  = 9'b111000010;
    mem[277]  = 9'b111000010;
    mem[278]  = 9'b111000010;
    mem[279]  = 9'b111000011;
    mem[280]  = 9'b111000011;
    mem[281]  = 9'b111000011;
    mem[282]  = 9'b111000011;
    mem[283]  = 9'b111000011;
    mem[284]  = 9'b111000100;
    mem[285]  = 9'b111000100;
    mem[286]  = 9'b111000100;
    mem[287]  = 9'b111000101;
    mem[288]  = 9'b111000101;
    mem[289]  = 9'b111000101;
    mem[290]  = 9'b111000101;
    mem[291]  = 9'b111000110;
    mem[292]  = 9'b111000110;
    mem[293]  = 9'b111000110;
    mem[294]  = 9'b111000111;
    mem[295]  = 9'b111000111;
    mem[296]  = 9'b111001000;
    mem[297]  = 9'b111001000;
    mem[298]  = 9'b111001000;
    mem[299]  = 9'b111001001;
    mem[300]  = 9'b111001001;
    mem[301]  = 9'b111001010;
    mem[302]  = 9'b111001010;
    mem[303]  = 9'b111001010;
    mem[304]  = 9'b111001011;
    mem[305]  = 9'b111001011;
    mem[306]  = 9'b111001100;
    mem[307]  = 9'b111001100;
    mem[308]  = 9'b111001101;
    mem[309]  = 9'b111001101;
    mem[310]  = 9'b111001110;
    mem[311]  = 9'b111001110;
    mem[312]  = 9'b111001111;
    mem[313]  = 9'b111001111;
    mem[314]  = 9'b111010000;
    mem[315]  = 9'b111010000;
    mem[316]  = 9'b111010001;
    mem[317]  = 9'b111010001;
    mem[318]  = 9'b111010010;
    mem[319]  = 9'b111010010;
    mem[320]  = 9'b111010011;
    mem[321]  = 9'b111010011;
    mem[322]  = 9'b111010100;
    mem[323]  = 9'b111010100;
    mem[324]  = 9'b111010101;
    mem[325]  = 9'b111010110;
    mem[326]  = 9'b111010110;
    mem[327]  = 9'b111010111;
    mem[328]  = 9'b111010111;
    mem[329]  = 9'b111011000;
    mem[330]  = 9'b111011001;
    mem[331]  = 9'b111011001;
    mem[332]  = 9'b111011010;
    mem[333]  = 9'b111011011;
    mem[334]  = 9'b111011011;
    mem[335]  = 9'b111011100;
    mem[336]  = 9'b111011100;
    mem[337]  = 9'b111011101;
    mem[338]  = 9'b111011110;
    mem[339]  = 9'b111011110;
    mem[340]  = 9'b111011111;
    mem[341]  = 9'b111100000;
    mem[342]  = 9'b111100000;
    mem[343]  = 9'b111100001;
    mem[344]  = 9'b111100010;
    mem[345]  = 9'b111100011;
    mem[346]  = 9'b111100011;
    mem[347]  = 9'b111100100;
    mem[348]  = 9'b111100101;
    mem[349]  = 9'b111100101;
    mem[350]  = 9'b111100110;
    mem[351]  = 9'b111100111;
    mem[352]  = 9'b111101000;
    mem[353]  = 9'b111101000;
    mem[354]  = 9'b111101001;
    mem[355]  = 9'b111101010;
    mem[356]  = 9'b111101010;
    mem[357]  = 9'b111101011;
    mem[358]  = 9'b111101100;
    mem[359]  = 9'b111101101;
    mem[360]  = 9'b111101101;
    mem[361]  = 9'b111101110;
    mem[362]  = 9'b111101111;
    mem[363]  = 9'b111110000;
    mem[364]  = 9'b111110000;
    mem[365]  = 9'b111110001;
    mem[366]  = 9'b111110010;
    mem[367]  = 9'b111110011;
    mem[368]  = 9'b111110100;
    mem[369]  = 9'b111110100;
    mem[370]  = 9'b111110101;
    mem[371]  = 9'b111110110;
    mem[372]  = 9'b111110111;
    mem[373]  = 9'b111110111;
    mem[374]  = 9'b111111000;
    mem[375]  = 9'b111111001;
    mem[376]  = 9'b111111010;
    mem[377]  = 9'b111111011;
    mem[378]  = 9'b111111011;
    mem[379]  = 9'b111111100;
    mem[380]  = 9'b111111101;
    mem[381]  = 9'b111111110;
    mem[382]  = 9'b111111110;
    mem[383]  = 9'b111111111;
    mem[384]  = 9'b000000000;
    mem[385]  = 9'b000000001;
    mem[386]  = 9'b000000010;
    mem[387]  = 9'b000000010;
    mem[388]  = 9'b000000011;
    mem[389]  = 9'b000000100;
    mem[390]  = 9'b000000101;
    mem[391]  = 9'b000000101;
    mem[392]  = 9'b000000110;
    mem[393]  = 9'b000000111;
    mem[394]  = 9'b000001000;
    mem[395]  = 9'b000001001;
    mem[396]  = 9'b000001001;
    mem[397]  = 9'b000001010;
    mem[398]  = 9'b000001011;
    mem[399]  = 9'b000001100;
    mem[400]  = 9'b000001100;
    mem[401]  = 9'b000001101;
    mem[402]  = 9'b000001110;
    mem[403]  = 9'b000001111;
    mem[404]  = 9'b000010000;
    mem[405]  = 9'b000010000;
    mem[406]  = 9'b000010001;
    mem[407]  = 9'b000010010;
    mem[408]  = 9'b000010011;
    mem[409]  = 9'b000010011;
    mem[410]  = 9'b000010100;
    mem[411]  = 9'b000010101;
    mem[412]  = 9'b000010110;
    mem[413]  = 9'b000010110;
    mem[414]  = 9'b000010111;
    mem[415]  = 9'b000011000;
    mem[416]  = 9'b000011000;
    mem[417]  = 9'b000011001;
    mem[418]  = 9'b000011010;
    mem[419]  = 9'b000011011;
    mem[420]  = 9'b000011011;
    mem[421]  = 9'b000011100;
    mem[422]  = 9'b000011101;
    mem[423]  = 9'b000011101;
    mem[424]  = 9'b000011110;
    mem[425]  = 9'b000011111;
    mem[426]  = 9'b000100000;
    mem[427]  = 9'b000100000;
    mem[428]  = 9'b000100001;
    mem[429]  = 9'b000100010;
    mem[430]  = 9'b000100010;
    mem[431]  = 9'b000100011;
    mem[432]  = 9'b000100100;
    mem[433]  = 9'b000100100;
    mem[434]  = 9'b000100101;
    mem[435]  = 9'b000100101;
    mem[436]  = 9'b000100110;
    mem[437]  = 9'b000100111;
    mem[438]  = 9'b000100111;
    mem[439]  = 9'b000101000;
    mem[440]  = 9'b000101001;
    mem[441]  = 9'b000101001;
    mem[442]  = 9'b000101010;
    mem[443]  = 9'b000101010;
    mem[444]  = 9'b000101011;
    mem[445]  = 9'b000101100;
    mem[446]  = 9'b000101100;
    mem[447]  = 9'b000101101;
    mem[448]  = 9'b000101101;
    mem[449]  = 9'b000101110;
    mem[450]  = 9'b000101110;
    mem[451]  = 9'b000101111;
    mem[452]  = 9'b000101111;
    mem[453]  = 9'b000110000;
    mem[454]  = 9'b000110000;
    mem[455]  = 9'b000110001;
    mem[456]  = 9'b000110001;
    mem[457]  = 9'b000110010;
    mem[458]  = 9'b000110010;
    mem[459]  = 9'b000110011;
    mem[460]  = 9'b000110011;
    mem[461]  = 9'b000110100;
    mem[462]  = 9'b000110100;
    mem[463]  = 9'b000110101;
    mem[464]  = 9'b000110101;
    mem[465]  = 9'b000110110;
    mem[466]  = 9'b000110110;
    mem[467]  = 9'b000110110;
    mem[468]  = 9'b000110111;
    mem[469]  = 9'b000110111;
    mem[470]  = 9'b000111000;
    mem[471]  = 9'b000111000;
    mem[472]  = 9'b000111000;
    mem[473]  = 9'b000111001;
    mem[474]  = 9'b000111001;
    mem[475]  = 9'b000111010;
    mem[476]  = 9'b000111010;
    mem[477]  = 9'b000111010;
    mem[478]  = 9'b000111011;
    mem[479]  = 9'b000111011;
    mem[480]  = 9'b000111011;
    mem[481]  = 9'b000111011;
    mem[482]  = 9'b000111100;
    mem[483]  = 9'b000111100;
    mem[484]  = 9'b000111100;
    mem[485]  = 9'b000111101;
    mem[486]  = 9'b000111101;
    mem[487]  = 9'b000111101;
    mem[488]  = 9'b000111101;
    mem[489]  = 9'b000111101;
    mem[490]  = 9'b000111110;
    mem[491]  = 9'b000111110;
    mem[492]  = 9'b000111110;
    mem[493]  = 9'b000111110;
    mem[494]  = 9'b000111110;
    mem[495]  = 9'b000111111;
    mem[496]  = 9'b000111111;
    mem[497]  = 9'b000111111;
    mem[498]  = 9'b000111111;
    mem[499]  = 9'b000111111;
    mem[500]  = 9'b000111111;
    mem[501]  = 9'b000111111;
    mem[502]  = 9'b001000000;
    mem[503]  = 9'b001000000;
    mem[504]  = 9'b001000000;
    mem[505]  = 9'b001000000;
    mem[506]  = 9'b001000000;
    mem[507]  = 9'b001000000;
    mem[508]  = 9'b001000000;
    mem[509]  = 9'b001000000;
    mem[510]  = 9'b001000000;
    mem[511]  = 9'b001000000;
  end

  // 동기식 출력
always_ff @(posedge clk) begin
  data[0]  <= mem[addr + 0];
  data[1]  <= mem[addr + 1];
  data[2]  <= mem[addr + 2];
  data[3]  <= mem[addr + 3];
  data[4]  <= mem[addr + 4];
  data[5]  <= mem[addr + 5];
  data[6]  <= mem[addr + 6];
  data[7]  <= mem[addr + 7];
  data[8]  <= mem[addr + 8];
  data[9]  <= mem[addr + 9];
  data[10] <= mem[addr + 10];
  data[11] <= mem[addr + 11];
  data[12] <= mem[addr + 12];
  data[13] <= mem[addr + 13];
  data[14] <= mem[addr + 14];
  data[15] <= mem[addr + 15];
end


endmodule

