`timescale 1ns/1ps

module twf_0_rom (
    input  logic         clk,
    input  logic         rstn,
    input  logic  [8:0]  address,           // base address
    output logic signed [8:0] twf_re[0:15], // 16개의 twiddle real
    output logic signed [8:0] twf_im[0:15]  // 16개의 twiddle imag
);

    // Twiddle factor ROM
    logic signed [8:0] twf_m0_re[0:511];
    logic signed [8:0] twf_m0_im[0:511];

    integer i;

    always_ff @(posedge clk or negedge rstn) begin
        if (!rstn) begin
            for (i = 0; i < 16; i++) begin
                twf_re[i] <= '0;
                twf_im[i] <= '0;
            end
        end else begin
            for (i = 0; i < 16; i++) begin
                twf_re[i] <= twf_m0_re[address + i];
                twf_im[i] <= twf_m0_im[address + i];
            end
        end
    end

    assign twf_m0_re[  0] = 128;    assign twf_m0_im[0] = 0;
    assign twf_m0_re[  1] = 128;    assign twf_m0_im[1] = 0;
    assign twf_m0_re[  2] = 128;    assign twf_m0_im[2] = 0;
    assign twf_m0_re[  3] = 128;    assign twf_m0_im[3] = 0;
    assign twf_m0_re[  4] = 128;    assign twf_m0_im[4] = 0;
    assign twf_m0_re[  5] = 128;    assign twf_m0_im[5] = 0;
    assign twf_m0_re[  6] = 128;    assign twf_m0_im[6] = 0;
    assign twf_m0_re[  7] = 128;    assign twf_m0_im[7] = 0;
    assign twf_m0_re[  8] = 128;    assign twf_m0_im[8] = 0;
    assign twf_m0_re[  9] = 128;    assign twf_m0_im[9] = 0;
    assign twf_m0_re[ 10] = 128;    assign twf_m0_im[10] = 0;
    assign twf_m0_re[ 11] = 128;    assign twf_m0_im[11] = 0;
    assign twf_m0_re[ 12] = 128;    assign twf_m0_im[12] = 0;
    assign twf_m0_re[ 13] = 128;    assign twf_m0_im[13] = 0;
    assign twf_m0_re[ 14] = 128;    assign twf_m0_im[14] = 0;
    assign twf_m0_re[ 15] = 128;    assign twf_m0_im[15] = 0;
    assign twf_m0_re[ 16] = 128;    assign twf_m0_im[16] = 0;
    assign twf_m0_re[ 17] = 128;    assign twf_m0_im[17] = 0;
    assign twf_m0_re[ 18] = 128;    assign twf_m0_im[18] = 0;
    assign twf_m0_re[ 19] = 128;    assign twf_m0_im[19] = 0;
    assign twf_m0_re[ 20] = 128;    assign twf_m0_im[20] = 0;
    assign twf_m0_re[ 21] = 128;    assign twf_m0_im[21] = 0;
    assign twf_m0_re[ 22] = 128;    assign twf_m0_im[22] = 0;
    assign twf_m0_re[ 23] = 128;    assign twf_m0_im[23] = 0;
    assign twf_m0_re[ 24] = 128;    assign twf_m0_im[24] = 0;
    assign twf_m0_re[ 25] = 128;    assign twf_m0_im[25] = 0;
    assign twf_m0_re[ 26] = 128;    assign twf_m0_im[26] = 0;
    assign twf_m0_re[ 27] = 128;    assign twf_m0_im[27] = 0;
    assign twf_m0_re[ 28] = 128;    assign twf_m0_im[28] = 0;
    assign twf_m0_re[ 29] = 128;    assign twf_m0_im[29] = 0;
    assign twf_m0_re[ 30] = 128;    assign twf_m0_im[30] = 0;
    assign twf_m0_re[ 31] = 128;    assign twf_m0_im[31] = 0;
    assign twf_m0_re[ 32] = 128;    assign twf_m0_im[32] = 0;
    assign twf_m0_re[ 33] = 128;    assign twf_m0_im[33] = 0;
    assign twf_m0_re[ 34] = 128;    assign twf_m0_im[34] = 0;
    assign twf_m0_re[ 35] = 128;    assign twf_m0_im[35] = 0;
    assign twf_m0_re[ 36] = 128;    assign twf_m0_im[36] = 0;
    assign twf_m0_re[ 37] = 128;    assign twf_m0_im[37] = 0;
    assign twf_m0_re[ 38] = 128;    assign twf_m0_im[38] = 0;
    assign twf_m0_re[ 39] = 128;    assign twf_m0_im[39] = 0;
    assign twf_m0_re[ 40] = 128;    assign twf_m0_im[40] = 0;
    assign twf_m0_re[ 41] = 128;    assign twf_m0_im[41] = 0;
    assign twf_m0_re[ 42] = 128;    assign twf_m0_im[42] = 0;
    assign twf_m0_re[ 43] = 128;    assign twf_m0_im[43] = 0;
    assign twf_m0_re[ 44] = 128;    assign twf_m0_im[44] = 0;
    assign twf_m0_re[ 45] = 128;    assign twf_m0_im[45] = 0;
    assign twf_m0_re[ 46] = 128;    assign twf_m0_im[46] = 0;
    assign twf_m0_re[ 47] = 128;    assign twf_m0_im[47] = 0;
    assign twf_m0_re[ 48] = 128;    assign twf_m0_im[48] = 0;
    assign twf_m0_re[ 49] = 128;    assign twf_m0_im[49] = 0;
    assign twf_m0_re[ 50] = 128;    assign twf_m0_im[50] = 0;
    assign twf_m0_re[ 51] = 128;    assign twf_m0_im[51] = 0;
    assign twf_m0_re[ 52] = 128;    assign twf_m0_im[52] = 0;
    assign twf_m0_re[ 53] = 128;    assign twf_m0_im[53] = 0;
    assign twf_m0_re[ 54] = 128;    assign twf_m0_im[54] = 0;
    assign twf_m0_re[ 55] = 128;    assign twf_m0_im[55] = 0;
    assign twf_m0_re[ 56] = 128;    assign twf_m0_im[56] = 0;
    assign twf_m0_re[ 57] = 128;    assign twf_m0_im[57] = 0;
    assign twf_m0_re[ 58] = 128;    assign twf_m0_im[58] = 0;
    assign twf_m0_re[ 59] = 128;    assign twf_m0_im[59] = 0;
    assign twf_m0_re[ 60] = 128;    assign twf_m0_im[60] = 0;
    assign twf_m0_re[ 61] = 128;    assign twf_m0_im[61] = 0;
    assign twf_m0_re[ 62] = 128;    assign twf_m0_im[62] = 0;
    assign twf_m0_re[ 63] = 128;    assign twf_m0_im[63] = 0;
    assign twf_m0_re[ 64] = 128;    assign twf_m0_im[64] = 0;
    assign twf_m0_re[ 65] = 128;    assign twf_m0_im[65] = -6;
    assign twf_m0_re[ 66] = 127;    assign twf_m0_im[66] = -13;
    assign twf_m0_re[ 67] = 127;    assign twf_m0_im[67] = -19;
    assign twf_m0_re[ 68] = 126;    assign twf_m0_im[68] = -25;
    assign twf_m0_re[ 69] = 124;    assign twf_m0_im[69] = -31;
    assign twf_m0_re[ 70] = 122;    assign twf_m0_im[70] = -37;
    assign twf_m0_re[ 71] = 121;    assign twf_m0_im[71] = -43;
    assign twf_m0_re[ 72] = 118;    assign twf_m0_im[72] = -49;
    assign twf_m0_re[ 73] = 116;    assign twf_m0_im[73] = -55;
    assign twf_m0_re[ 74] = 113;    assign twf_m0_im[74] = -60;
    assign twf_m0_re[ 75] = 110;    assign twf_m0_im[75] = -66;
    assign twf_m0_re[ 76] = 106;    assign twf_m0_im[76] = -71;
    assign twf_m0_re[ 77] = 103;    assign twf_m0_im[77] = -76;
    assign twf_m0_re[ 78] = 99;    assign twf_m0_im[78] = -81;
    assign twf_m0_re[ 79] = 95;    assign twf_m0_im[79] = -86;
    assign twf_m0_re[ 80] = 91;    assign twf_m0_im[80] = -91;
    assign twf_m0_re[ 81] = 86;    assign twf_m0_im[81] = -95;
    assign twf_m0_re[ 82] = 81;    assign twf_m0_im[82] = -99;
    assign twf_m0_re[ 83] = 76;    assign twf_m0_im[83] = -103;
    assign twf_m0_re[ 84] = 71;    assign twf_m0_im[84] = -106;
    assign twf_m0_re[ 85] = 66;    assign twf_m0_im[85] = -110;
    assign twf_m0_re[ 86] = 60;    assign twf_m0_im[86] = -113;
    assign twf_m0_re[ 87] = 55;    assign twf_m0_im[87] = -116;
    assign twf_m0_re[ 88] = 49;    assign twf_m0_im[88] = -118;
    assign twf_m0_re[ 89] = 43;    assign twf_m0_im[89] = -121;
    assign twf_m0_re[ 90] = 37;    assign twf_m0_im[90] = -122;
    assign twf_m0_re[ 91] = 31;    assign twf_m0_im[91] = -124;
    assign twf_m0_re[ 92] = 25;    assign twf_m0_im[92] = -126;
    assign twf_m0_re[ 93] = 19;    assign twf_m0_im[93] = -127;
    assign twf_m0_re[ 94] = 13;    assign twf_m0_im[94] = -127;
    assign twf_m0_re[ 95] = 6;    assign twf_m0_im[95] = -128;
    assign twf_m0_re[ 96] = 0;    assign twf_m0_im[96] = -128;
    assign twf_m0_re[ 97] = -6;    assign twf_m0_im[97] = -128;
    assign twf_m0_re[ 98] = -13;    assign twf_m0_im[98] = -127;
    assign twf_m0_re[ 99] = -19;    assign twf_m0_im[99] = -127;
    assign twf_m0_re[100] = -25;    assign twf_m0_im[100] = -126;
    assign twf_m0_re[101] = -31;    assign twf_m0_im[101] = -124;
    assign twf_m0_re[102] = -37;    assign twf_m0_im[102] = -122;
    assign twf_m0_re[103] = -43;    assign twf_m0_im[103] = -121;
    assign twf_m0_re[104] = -49;    assign twf_m0_im[104] = -118;
    assign twf_m0_re[105] = -55;    assign twf_m0_im[105] = -116;
    assign twf_m0_re[106] = -60;    assign twf_m0_im[106] = -113;
    assign twf_m0_re[107] = -66;    assign twf_m0_im[107] = -110;
    assign twf_m0_re[108] = -71;    assign twf_m0_im[108] = -106;
    assign twf_m0_re[109] = -76;    assign twf_m0_im[109] = -103;
    assign twf_m0_re[110] = -81;    assign twf_m0_im[110] = -99;
    assign twf_m0_re[111] = -86;    assign twf_m0_im[111] = -95;
    assign twf_m0_re[112] = -91;    assign twf_m0_im[112] = -91;
    assign twf_m0_re[113] = -95;    assign twf_m0_im[113] = -86;
    assign twf_m0_re[114] = -99;    assign twf_m0_im[114] = -81;
    assign twf_m0_re[115] = -103;    assign twf_m0_im[115] = -76;
    assign twf_m0_re[116] = -106;    assign twf_m0_im[116] = -71;
    assign twf_m0_re[117] = -110;    assign twf_m0_im[117] = -66;
    assign twf_m0_re[118] = -113;    assign twf_m0_im[118] = -60;
    assign twf_m0_re[119] = -116;    assign twf_m0_im[119] = -55;
    assign twf_m0_re[120] = -118;    assign twf_m0_im[120] = -49;
    assign twf_m0_re[121] = -121;    assign twf_m0_im[121] = -43;
    assign twf_m0_re[122] = -122;    assign twf_m0_im[122] = -37;
    assign twf_m0_re[123] = -124;    assign twf_m0_im[123] = -31;
    assign twf_m0_re[124] = -126;    assign twf_m0_im[124] = -25;
    assign twf_m0_re[125] = -127;    assign twf_m0_im[125] = -19;
    assign twf_m0_re[126] = -127;    assign twf_m0_im[126] = -13;
    assign twf_m0_re[127] = -128;    assign twf_m0_im[127] = -6;
    assign twf_m0_re[128] = 128;    assign twf_m0_im[128] = 0;
    assign twf_m0_re[129] = 128;    assign twf_m0_im[129] = -3;
    assign twf_m0_re[130] = 128;    assign twf_m0_im[130] = -6;
    assign twf_m0_re[131] = 128;    assign twf_m0_im[131] = -9;
    assign twf_m0_re[132] = 127;    assign twf_m0_im[132] = -13;
    assign twf_m0_re[133] = 127;    assign twf_m0_im[133] = -16;
    assign twf_m0_re[134] = 127;    assign twf_m0_im[134] = -19;
    assign twf_m0_re[135] = 126;    assign twf_m0_im[135] = -22;
    assign twf_m0_re[136] = 126;    assign twf_m0_im[136] = -25;
    assign twf_m0_re[137] = 125;    assign twf_m0_im[137] = -28;
    assign twf_m0_re[138] = 124;    assign twf_m0_im[138] = -31;
    assign twf_m0_re[139] = 123;    assign twf_m0_im[139] = -34;
    assign twf_m0_re[140] = 122;    assign twf_m0_im[140] = -37;
    assign twf_m0_re[141] = 122;    assign twf_m0_im[141] = -40;
    assign twf_m0_re[142] = 121;    assign twf_m0_im[142] = -43;
    assign twf_m0_re[143] = 119;    assign twf_m0_im[143] = -46;
    assign twf_m0_re[144] = 118;    assign twf_m0_im[144] = -49;
    assign twf_m0_re[145] = 117;    assign twf_m0_im[145] = -52;
    assign twf_m0_re[146] = 116;    assign twf_m0_im[146] = -55;
    assign twf_m0_re[147] = 114;    assign twf_m0_im[147] = -58;
    assign twf_m0_re[148] = 113;    assign twf_m0_im[148] = -60;
    assign twf_m0_re[149] = 111;    assign twf_m0_im[149] = -63;
    assign twf_m0_re[150] = 110;    assign twf_m0_im[150] = -66;
    assign twf_m0_re[151] = 108;    assign twf_m0_im[151] = -68;
    assign twf_m0_re[152] = 106;    assign twf_m0_im[152] = -71;
    assign twf_m0_re[153] = 105;    assign twf_m0_im[153] = -74;
    assign twf_m0_re[154] = 103;    assign twf_m0_im[154] = -76;
    assign twf_m0_re[155] = 101;    assign twf_m0_im[155] = -79;
    assign twf_m0_re[156] = 99;    assign twf_m0_im[156] = -81;
    assign twf_m0_re[157] = 97;    assign twf_m0_im[157] = -84;
    assign twf_m0_re[158] = 95;    assign twf_m0_im[158] = -86;
    assign twf_m0_re[159] = 93;    assign twf_m0_im[159] = -88;
    assign twf_m0_re[160] = 91;    assign twf_m0_im[160] = -91;
    assign twf_m0_re[161] = 88;    assign twf_m0_im[161] = -93;
    assign twf_m0_re[162] = 86;    assign twf_m0_im[162] = -95;
    assign twf_m0_re[163] = 84;    assign twf_m0_im[163] = -97;
    assign twf_m0_re[164] = 81;    assign twf_m0_im[164] = -99;
    assign twf_m0_re[165] = 79;    assign twf_m0_im[165] = -101;
    assign twf_m0_re[166] = 76;    assign twf_m0_im[166] = -103;
    assign twf_m0_re[167] = 74;    assign twf_m0_im[167] = -105;
    assign twf_m0_re[168] = 71;    assign twf_m0_im[168] = -106;
    assign twf_m0_re[169] = 68;    assign twf_m0_im[169] = -108;
    assign twf_m0_re[170] = 66;    assign twf_m0_im[170] = -110;
    assign twf_m0_re[171] = 63;    assign twf_m0_im[171] = -111;
    assign twf_m0_re[172] = 60;    assign twf_m0_im[172] = -113;
    assign twf_m0_re[173] = 58;    assign twf_m0_im[173] = -114;
    assign twf_m0_re[174] = 55;    assign twf_m0_im[174] = -116;
    assign twf_m0_re[175] = 52;    assign twf_m0_im[175] = -117;
    assign twf_m0_re[176] = 49;    assign twf_m0_im[176] = -118;
    assign twf_m0_re[177] = 46;    assign twf_m0_im[177] = -119;
    assign twf_m0_re[178] = 43;    assign twf_m0_im[178] = -121;
    assign twf_m0_re[179] = 40;    assign twf_m0_im[179] = -122;
    assign twf_m0_re[180] = 37;    assign twf_m0_im[180] = -122;
    assign twf_m0_re[181] = 34;    assign twf_m0_im[181] = -123;
    assign twf_m0_re[182] = 31;    assign twf_m0_im[182] = -124;
    assign twf_m0_re[183] = 28;    assign twf_m0_im[183] = -125;
    assign twf_m0_re[184] = 25;    assign twf_m0_im[184] = -126;
    assign twf_m0_re[185] = 22;    assign twf_m0_im[185] = -126;
    assign twf_m0_re[186] = 19;    assign twf_m0_im[186] = -127;
    assign twf_m0_re[187] = 16;    assign twf_m0_im[187] = -127;
    assign twf_m0_re[188] = 13;    assign twf_m0_im[188] = -127;
    assign twf_m0_re[189] = 9;    assign twf_m0_im[189] = -128;
    assign twf_m0_re[190] = 6;    assign twf_m0_im[190] = -128;
    assign twf_m0_re[191] = 3;    assign twf_m0_im[191] = -128;
    assign twf_m0_re[192] = 128;    assign twf_m0_im[192] = 0;
    assign twf_m0_re[193] = 128;    assign twf_m0_im[193] = -9;
    assign twf_m0_re[194] = 127;    assign twf_m0_im[194] = -19;
    assign twf_m0_re[195] = 125;    assign twf_m0_im[195] = -28;
    assign twf_m0_re[196] = 122;    assign twf_m0_im[196] = -37;
    assign twf_m0_re[197] = 119;    assign twf_m0_im[197] = -46;
    assign twf_m0_re[198] = 116;    assign twf_m0_im[198] = -55;
    assign twf_m0_re[199] = 111;    assign twf_m0_im[199] = -63;
    assign twf_m0_re[200] = 106;    assign twf_m0_im[200] = -71;
    assign twf_m0_re[201] = 101;    assign twf_m0_im[201] = -79;
    assign twf_m0_re[202] = 95;    assign twf_m0_im[202] = -86;
    assign twf_m0_re[203] = 88;    assign twf_m0_im[203] = -93;
    assign twf_m0_re[204] = 81;    assign twf_m0_im[204] = -99;
    assign twf_m0_re[205] = 74;    assign twf_m0_im[205] = -105;
    assign twf_m0_re[206] = 66;    assign twf_m0_im[206] = -110;
    assign twf_m0_re[207] = 58;    assign twf_m0_im[207] = -114;
    assign twf_m0_re[208] = 49;    assign twf_m0_im[208] = -118;
    assign twf_m0_re[209] = 40;    assign twf_m0_im[209] = -122;
    assign twf_m0_re[210] = 31;    assign twf_m0_im[210] = -124;
    assign twf_m0_re[211] = 22;    assign twf_m0_im[211] = -126;
    assign twf_m0_re[212] = 13;    assign twf_m0_im[212] = -127;
    assign twf_m0_re[213] = 3;    assign twf_m0_im[213] = -128;
    assign twf_m0_re[214] = -6;    assign twf_m0_im[214] = -128;
    assign twf_m0_re[215] = -16;    assign twf_m0_im[215] = -127;
    assign twf_m0_re[216] = -25;    assign twf_m0_im[216] = -126;
    assign twf_m0_re[217] = -34;    assign twf_m0_im[217] = -123;
    assign twf_m0_re[218] = -43;    assign twf_m0_im[218] = -121;
    assign twf_m0_re[219] = -52;    assign twf_m0_im[219] = -117;
    assign twf_m0_re[220] = -60;    assign twf_m0_im[220] = -113;
    assign twf_m0_re[221] = -68;    assign twf_m0_im[221] = -108;
    assign twf_m0_re[222] = -76;    assign twf_m0_im[222] = -103;
    assign twf_m0_re[223] = -84;    assign twf_m0_im[223] = -97;
    assign twf_m0_re[224] = -91;    assign twf_m0_im[224] = -91;
    assign twf_m0_re[225] = -97;    assign twf_m0_im[225] = -84;
    assign twf_m0_re[226] = -103;    assign twf_m0_im[226] = -76;
    assign twf_m0_re[227] = -108;    assign twf_m0_im[227] = -68;
    assign twf_m0_re[228] = -113;    assign twf_m0_im[228] = -60;
    assign twf_m0_re[229] = -117;    assign twf_m0_im[229] = -52;
    assign twf_m0_re[230] = -121;    assign twf_m0_im[230] = -43;
    assign twf_m0_re[231] = -123;    assign twf_m0_im[231] = -34;
    assign twf_m0_re[232] = -126;    assign twf_m0_im[232] = -25;
    assign twf_m0_re[233] = -127;    assign twf_m0_im[233] = -16;
    assign twf_m0_re[234] = -128;    assign twf_m0_im[234] = -6;
    assign twf_m0_re[235] = -128;    assign twf_m0_im[235] = 3;
    assign twf_m0_re[236] = -127;    assign twf_m0_im[236] = 13;
    assign twf_m0_re[237] = -126;    assign twf_m0_im[237] = 22;
    assign twf_m0_re[238] = -124;    assign twf_m0_im[238] = 31;
    assign twf_m0_re[239] = -122;    assign twf_m0_im[239] = 40;
    assign twf_m0_re[240] = -118;    assign twf_m0_im[240] = 49;
    assign twf_m0_re[241] = -114;    assign twf_m0_im[241] = 58;
    assign twf_m0_re[242] = -110;    assign twf_m0_im[242] = 66;
    assign twf_m0_re[243] = -105;    assign twf_m0_im[243] = 74;
    assign twf_m0_re[244] = -99;    assign twf_m0_im[244] = 81;
    assign twf_m0_re[245] = -93;    assign twf_m0_im[245] = 88;
    assign twf_m0_re[246] = -86;    assign twf_m0_im[246] = 95;
    assign twf_m0_re[247] = -79;    assign twf_m0_im[247] = 101;
    assign twf_m0_re[248] = -71;    assign twf_m0_im[248] = 106;
    assign twf_m0_re[249] = -63;    assign twf_m0_im[249] = 111;
    assign twf_m0_re[250] = -55;    assign twf_m0_im[250] = 116;
    assign twf_m0_re[251] = -46;    assign twf_m0_im[251] = 119;
    assign twf_m0_re[252] = -37;    assign twf_m0_im[252] = 122;
    assign twf_m0_re[253] = -28;    assign twf_m0_im[253] = 125;
    assign twf_m0_re[254] = -19;    assign twf_m0_im[254] = 127;
    assign twf_m0_re[255] = -9;    assign twf_m0_im[255] = 128;
    assign twf_m0_re[256] = 128;    assign twf_m0_im[256] = 0;
    assign twf_m0_re[257] = 128;    assign twf_m0_im[257] = -2;
    assign twf_m0_re[258] = 128;    assign twf_m0_im[258] = -3;
    assign twf_m0_re[259] = 128;    assign twf_m0_im[259] = -5;
    assign twf_m0_re[260] = 128;    assign twf_m0_im[260] = -6;
    assign twf_m0_re[261] = 128;    assign twf_m0_im[261] = -8;
    assign twf_m0_re[262] = 128;    assign twf_m0_im[262] = -9;
    assign twf_m0_re[263] = 128;    assign twf_m0_im[263] = -11;
    assign twf_m0_re[264] = 127;    assign twf_m0_im[264] = -13;
    assign twf_m0_re[265] = 127;    assign twf_m0_im[265] = -14;
    assign twf_m0_re[266] = 127;    assign twf_m0_im[266] = -16;
    assign twf_m0_re[267] = 127;    assign twf_m0_im[267] = -17;
    assign twf_m0_re[268] = 127;    assign twf_m0_im[268] = -19;
    assign twf_m0_re[269] = 126;    assign twf_m0_im[269] = -20;
    assign twf_m0_re[270] = 126;    assign twf_m0_im[270] = -22;
    assign twf_m0_re[271] = 126;    assign twf_m0_im[271] = -23;
    assign twf_m0_re[272] = 126;    assign twf_m0_im[272] = -25;
    assign twf_m0_re[273] = 125;    assign twf_m0_im[273] = -27;
    assign twf_m0_re[274] = 125;    assign twf_m0_im[274] = -28;
    assign twf_m0_re[275] = 125;    assign twf_m0_im[275] = -30;
    assign twf_m0_re[276] = 124;    assign twf_m0_im[276] = -31;
    assign twf_m0_re[277] = 124;    assign twf_m0_im[277] = -33;
    assign twf_m0_re[278] = 123;    assign twf_m0_im[278] = -34;
    assign twf_m0_re[279] = 123;    assign twf_m0_im[279] = -36;
    assign twf_m0_re[280] = 122;    assign twf_m0_im[280] = -37;
    assign twf_m0_re[281] = 122;    assign twf_m0_im[281] = -39;
    assign twf_m0_re[282] = 122;    assign twf_m0_im[282] = -40;
    assign twf_m0_re[283] = 121;    assign twf_m0_im[283] = -42;
    assign twf_m0_re[284] = 121;    assign twf_m0_im[284] = -43;
    assign twf_m0_re[285] = 120;    assign twf_m0_im[285] = -45;
    assign twf_m0_re[286] = 119;    assign twf_m0_im[286] = -46;
    assign twf_m0_re[287] = 119;    assign twf_m0_im[287] = -48;
    assign twf_m0_re[288] = 118;    assign twf_m0_im[288] = -49;
    assign twf_m0_re[289] = 118;    assign twf_m0_im[289] = -50;
    assign twf_m0_re[290] = 117;    assign twf_m0_im[290] = -52;
    assign twf_m0_re[291] = 116;    assign twf_m0_im[291] = -53;
    assign twf_m0_re[292] = 116;    assign twf_m0_im[292] = -55;
    assign twf_m0_re[293] = 115;    assign twf_m0_im[293] = -56;
    assign twf_m0_re[294] = 114;    assign twf_m0_im[294] = -58;
    assign twf_m0_re[295] = 114;    assign twf_m0_im[295] = -59;
    assign twf_m0_re[296] = 113;    assign twf_m0_im[296] = -60;
    assign twf_m0_re[297] = 112;    assign twf_m0_im[297] = -62;
    assign twf_m0_re[298] = 111;    assign twf_m0_im[298] = -63;
    assign twf_m0_re[299] = 111;    assign twf_m0_im[299] = -64;
    assign twf_m0_re[300] = 110;    assign twf_m0_im[300] = -66;
    assign twf_m0_re[301] = 109;    assign twf_m0_im[301] = -67;
    assign twf_m0_re[302] = 108;    assign twf_m0_im[302] = -68;
    assign twf_m0_re[303] = 107;    assign twf_m0_im[303] = -70;
    assign twf_m0_re[304] = 106;    assign twf_m0_im[304] = -71;
    assign twf_m0_re[305] = 106;    assign twf_m0_im[305] = -72;
    assign twf_m0_re[306] = 105;    assign twf_m0_im[306] = -74;
    assign twf_m0_re[307] = 104;    assign twf_m0_im[307] = -75;
    assign twf_m0_re[308] = 103;    assign twf_m0_im[308] = -76;
    assign twf_m0_re[309] = 102;    assign twf_m0_im[309] = -78;
    assign twf_m0_re[310] = 101;    assign twf_m0_im[310] = -79;
    assign twf_m0_re[311] = 100;    assign twf_m0_im[311] = -80;
    assign twf_m0_re[312] = 99;    assign twf_m0_im[312] = -81;
    assign twf_m0_re[313] = 98;    assign twf_m0_im[313] = -82;
    assign twf_m0_re[314] = 97;    assign twf_m0_im[314] = -84;
    assign twf_m0_re[315] = 96;    assign twf_m0_im[315] = -85;
    assign twf_m0_re[316] = 95;    assign twf_m0_im[316] = -86;
    assign twf_m0_re[317] = 94;    assign twf_m0_im[317] = -87;
    assign twf_m0_re[318] = 93;    assign twf_m0_im[318] = -88;
    assign twf_m0_re[319] = 92;    assign twf_m0_im[319] = -89;
    assign twf_m0_re[320] = 128;    assign twf_m0_im[320] = 0;
    assign twf_m0_re[321] = 128;    assign twf_m0_im[321] = -8;
    assign twf_m0_re[322] = 127;    assign twf_m0_im[322] = -16;
    assign twf_m0_re[323] = 126;    assign twf_m0_im[323] = -23;
    assign twf_m0_re[324] = 124;    assign twf_m0_im[324] = -31;
    assign twf_m0_re[325] = 122;    assign twf_m0_im[325] = -39;
    assign twf_m0_re[326] = 119;    assign twf_m0_im[326] = -46;
    assign twf_m0_re[327] = 116;    assign twf_m0_im[327] = -53;
    assign twf_m0_re[328] = 113;    assign twf_m0_im[328] = -60;
    assign twf_m0_re[329] = 109;    assign twf_m0_im[329] = -67;
    assign twf_m0_re[330] = 105;    assign twf_m0_im[330] = -74;
    assign twf_m0_re[331] = 100;    assign twf_m0_im[331] = -80;
    assign twf_m0_re[332] = 95;    assign twf_m0_im[332] = -86;
    assign twf_m0_re[333] = 89;    assign twf_m0_im[333] = -92;
    assign twf_m0_re[334] = 84;    assign twf_m0_im[334] = -97;
    assign twf_m0_re[335] = 78;    assign twf_m0_im[335] = -102;
    assign twf_m0_re[336] = 71;    assign twf_m0_im[336] = -106;
    assign twf_m0_re[337] = 64;    assign twf_m0_im[337] = -111;
    assign twf_m0_re[338] = 58;    assign twf_m0_im[338] = -114;
    assign twf_m0_re[339] = 50;    assign twf_m0_im[339] = -118;
    assign twf_m0_re[340] = 43;    assign twf_m0_im[340] = -121;
    assign twf_m0_re[341] = 36;    assign twf_m0_im[341] = -123;
    assign twf_m0_re[342] = 28;    assign twf_m0_im[342] = -125;
    assign twf_m0_re[343] = 20;    assign twf_m0_im[343] = -126;
    assign twf_m0_re[344] = 13;    assign twf_m0_im[344] = -127;
    assign twf_m0_re[345] = 5;    assign twf_m0_im[345] = -128;
    assign twf_m0_re[346] = -3;    assign twf_m0_im[346] = -128;
    assign twf_m0_re[347] = -11;    assign twf_m0_im[347] = -128;
    assign twf_m0_re[348] = -19;    assign twf_m0_im[348] = -127;
    assign twf_m0_re[349] = -27;    assign twf_m0_im[349] = -125;
    assign twf_m0_re[350] = -34;    assign twf_m0_im[350] = -123;
    assign twf_m0_re[351] = -42;    assign twf_m0_im[351] = -121;
    assign twf_m0_re[352] = -49;    assign twf_m0_im[352] = -118;
    assign twf_m0_re[353] = -56;    assign twf_m0_im[353] = -115;
    assign twf_m0_re[354] = -63;    assign twf_m0_im[354] = -111;
    assign twf_m0_re[355] = -70;    assign twf_m0_im[355] = -107;
    assign twf_m0_re[356] = -76;    assign twf_m0_im[356] = -103;
    assign twf_m0_re[357] = -82;    assign twf_m0_im[357] = -98;
    assign twf_m0_re[358] = -88;    assign twf_m0_im[358] = -93;
    assign twf_m0_re[359] = -94;    assign twf_m0_im[359] = -87;
    assign twf_m0_re[360] = -99;    assign twf_m0_im[360] = -81;
    assign twf_m0_re[361] = -104;    assign twf_m0_im[361] = -75;
    assign twf_m0_re[362] = -108;    assign twf_m0_im[362] = -68;
    assign twf_m0_re[363] = -112;    assign twf_m0_im[363] = -62;
    assign twf_m0_re[364] = -116;    assign twf_m0_im[364] = -55;
    assign twf_m0_re[365] = -119;    assign twf_m0_im[365] = -48;
    assign twf_m0_re[366] = -122;    assign twf_m0_im[366] = -40;
    assign twf_m0_re[367] = -124;    assign twf_m0_im[367] = -33;
    assign twf_m0_re[368] = -126;    assign twf_m0_im[368] = -25;
    assign twf_m0_re[369] = -127;    assign twf_m0_im[369] = -17;
    assign twf_m0_re[370] = -128;    assign twf_m0_im[370] = -9;
    assign twf_m0_re[371] = -128;    assign twf_m0_im[371] = -2;
    assign twf_m0_re[372] = -128;    assign twf_m0_im[372] = 6;
    assign twf_m0_re[373] = -127;    assign twf_m0_im[373] = 14;
    assign twf_m0_re[374] = -126;    assign twf_m0_im[374] = 22;
    assign twf_m0_re[375] = -125;    assign twf_m0_im[375] = 30;
    assign twf_m0_re[376] = -122;    assign twf_m0_im[376] = 37;
    assign twf_m0_re[377] = -120;    assign twf_m0_im[377] = 45;
    assign twf_m0_re[378] = -117;    assign twf_m0_im[378] = 52;
    assign twf_m0_re[379] = -114;    assign twf_m0_im[379] = 59;
    assign twf_m0_re[380] = -110;    assign twf_m0_im[380] = 66;
    assign twf_m0_re[381] = -106;    assign twf_m0_im[381] = 72;
    assign twf_m0_re[382] = -101;    assign twf_m0_im[382] = 79;
    assign twf_m0_re[383] = -96;    assign twf_m0_im[383] = 85;
    assign twf_m0_re[384] = 128;    assign twf_m0_im[384] = 0;
    assign twf_m0_re[385] = 128;    assign twf_m0_im[385] = -5;
    assign twf_m0_re[386] = 128;    assign twf_m0_im[386] = -9;
    assign twf_m0_re[387] = 127;    assign twf_m0_im[387] = -14;
    assign twf_m0_re[388] = 127;    assign twf_m0_im[388] = -19;
    assign twf_m0_re[389] = 126;    assign twf_m0_im[389] = -23;
    assign twf_m0_re[390] = 125;    assign twf_m0_im[390] = -28;
    assign twf_m0_re[391] = 124;    assign twf_m0_im[391] = -33;
    assign twf_m0_re[392] = 122;    assign twf_m0_im[392] = -37;
    assign twf_m0_re[393] = 121;    assign twf_m0_im[393] = -42;
    assign twf_m0_re[394] = 119;    assign twf_m0_im[394] = -46;
    assign twf_m0_re[395] = 118;    assign twf_m0_im[395] = -50;
    assign twf_m0_re[396] = 116;    assign twf_m0_im[396] = -55;
    assign twf_m0_re[397] = 114;    assign twf_m0_im[397] = -59;
    assign twf_m0_re[398] = 111;    assign twf_m0_im[398] = -63;
    assign twf_m0_re[399] = 109;    assign twf_m0_im[399] = -67;
    assign twf_m0_re[400] = 106;    assign twf_m0_im[400] = -71;
    assign twf_m0_re[401] = 104;    assign twf_m0_im[401] = -75;
    assign twf_m0_re[402] = 101;    assign twf_m0_im[402] = -79;
    assign twf_m0_re[403] = 98;    assign twf_m0_im[403] = -82;
    assign twf_m0_re[404] = 95;    assign twf_m0_im[404] = -86;
    assign twf_m0_re[405] = 92;    assign twf_m0_im[405] = -89;
    assign twf_m0_re[406] = 88;    assign twf_m0_im[406] = -93;
    assign twf_m0_re[407] = 85;    assign twf_m0_im[407] = -96;
    assign twf_m0_re[408] = 81;    assign twf_m0_im[408] = -99;
    assign twf_m0_re[409] = 78;    assign twf_m0_im[409] = -102;
    assign twf_m0_re[410] = 74;    assign twf_m0_im[410] = -105;
    assign twf_m0_re[411] = 70;    assign twf_m0_im[411] = -107;
    assign twf_m0_re[412] = 66;    assign twf_m0_im[412] = -110;
    assign twf_m0_re[413] = 62;    assign twf_m0_im[413] = -112;
    assign twf_m0_re[414] = 58;    assign twf_m0_im[414] = -114;
    assign twf_m0_re[415] = 53;    assign twf_m0_im[415] = -116;
    assign twf_m0_re[416] = 49;    assign twf_m0_im[416] = -118;
    assign twf_m0_re[417] = 45;    assign twf_m0_im[417] = -120;
    assign twf_m0_re[418] = 40;    assign twf_m0_im[418] = -122;
    assign twf_m0_re[419] = 36;    assign twf_m0_im[419] = -123;
    assign twf_m0_re[420] = 31;    assign twf_m0_im[420] = -124;
    assign twf_m0_re[421] = 27;    assign twf_m0_im[421] = -125;
    assign twf_m0_re[422] = 22;    assign twf_m0_im[422] = -126;
    assign twf_m0_re[423] = 17;    assign twf_m0_im[423] = -127;
    assign twf_m0_re[424] = 13;    assign twf_m0_im[424] = -127;
    assign twf_m0_re[425] = 8;    assign twf_m0_im[425] = -128;
    assign twf_m0_re[426] = 3;    assign twf_m0_im[426] = -128;
    assign twf_m0_re[427] = -2;    assign twf_m0_im[427] = -128;
    assign twf_m0_re[428] = -6;    assign twf_m0_im[428] = -128;
    assign twf_m0_re[429] = -11;    assign twf_m0_im[429] = -128;
    assign twf_m0_re[430] = -16;    assign twf_m0_im[430] = -127;
    assign twf_m0_re[431] = -20;    assign twf_m0_im[431] = -126;
    assign twf_m0_re[432] = -25;    assign twf_m0_im[432] = -126;
    assign twf_m0_re[433] = -30;    assign twf_m0_im[433] = -125;
    assign twf_m0_re[434] = -34;    assign twf_m0_im[434] = -123;
    assign twf_m0_re[435] = -39;    assign twf_m0_im[435] = -122;
    assign twf_m0_re[436] = -43;    assign twf_m0_im[436] = -121;
    assign twf_m0_re[437] = -48;    assign twf_m0_im[437] = -119;
    assign twf_m0_re[438] = -52;    assign twf_m0_im[438] = -117;
    assign twf_m0_re[439] = -56;    assign twf_m0_im[439] = -115;
    assign twf_m0_re[440] = -60;    assign twf_m0_im[440] = -113;
    assign twf_m0_re[441] = -64;    assign twf_m0_im[441] = -111;
    assign twf_m0_re[442] = -68;    assign twf_m0_im[442] = -108;
    assign twf_m0_re[443] = -72;    assign twf_m0_im[443] = -106;
    assign twf_m0_re[444] = -76;    assign twf_m0_im[444] = -103;
    assign twf_m0_re[445] = -80;    assign twf_m0_im[445] = -100;
    assign twf_m0_re[446] = -84;    assign twf_m0_im[446] = -97;
    assign twf_m0_re[447] = -87;    assign twf_m0_im[447] = -94;
    assign twf_m0_re[448] = 128;    assign twf_m0_im[448] = 0;
    assign twf_m0_re[449] = 128;    assign twf_m0_im[449] = -11;
    assign twf_m0_re[450] = 126;    assign twf_m0_im[450] = -22;
    assign twf_m0_re[451] = 124;    assign twf_m0_im[451] = -33;
    assign twf_m0_re[452] = 121;    assign twf_m0_im[452] = -43;
    assign twf_m0_re[453] = 116;    assign twf_m0_im[453] = -53;
    assign twf_m0_re[454] = 111;    assign twf_m0_im[454] = -63;
    assign twf_m0_re[455] = 106;    assign twf_m0_im[455] = -72;
    assign twf_m0_re[456] = 99;    assign twf_m0_im[456] = -81;
    assign twf_m0_re[457] = 92;    assign twf_m0_im[457] = -89;
    assign twf_m0_re[458] = 84;    assign twf_m0_im[458] = -97;
    assign twf_m0_re[459] = 75;    assign twf_m0_im[459] = -104;
    assign twf_m0_re[460] = 66;    assign twf_m0_im[460] = -110;
    assign twf_m0_re[461] = 56;    assign twf_m0_im[461] = -115;
    assign twf_m0_re[462] = 46;    assign twf_m0_im[462] = -119;
    assign twf_m0_re[463] = 36;    assign twf_m0_im[463] = -123;
    assign twf_m0_re[464] = 25;    assign twf_m0_im[464] = -126;
    assign twf_m0_re[465] = 14;    assign twf_m0_im[465] = -127;
    assign twf_m0_re[466] = 3;    assign twf_m0_im[466] = -128;
    assign twf_m0_re[467] = -8;    assign twf_m0_im[467] = -128;
    assign twf_m0_re[468] = -19;    assign twf_m0_im[468] = -127;
    assign twf_m0_re[469] = -30;    assign twf_m0_im[469] = -125;
    assign twf_m0_re[470] = -40;    assign twf_m0_im[470] = -122;
    assign twf_m0_re[471] = -50;    assign twf_m0_im[471] = -118;
    assign twf_m0_re[472] = -60;    assign twf_m0_im[472] = -113;
    assign twf_m0_re[473] = -70;    assign twf_m0_im[473] = -107;
    assign twf_m0_re[474] = -79;    assign twf_m0_im[474] = -101;
    assign twf_m0_re[475] = -87;    assign twf_m0_im[475] = -94;
    assign twf_m0_re[476] = -95;    assign twf_m0_im[476] = -86;
    assign twf_m0_re[477] = -102;    assign twf_m0_im[477] = -78;
    assign twf_m0_re[478] = -108;    assign twf_m0_im[478] = -68;
    assign twf_m0_re[479] = -114;    assign twf_m0_im[479] = -59;
    assign twf_m0_re[480] = -118;    assign twf_m0_im[480] = -49;
    assign twf_m0_re[481] = -122;    assign twf_m0_im[481] = -39;
    assign twf_m0_re[482] = -125;    assign twf_m0_im[482] = -28;
    assign twf_m0_re[483] = -127;    assign twf_m0_im[483] = -17;
    assign twf_m0_re[484] = -128;    assign twf_m0_im[484] = -6;
    assign twf_m0_re[485] = -128;    assign twf_m0_im[485] = 5;
    assign twf_m0_re[486] = -127;    assign twf_m0_im[486] = 16;
    assign twf_m0_re[487] = -125;    assign twf_m0_im[487] = 27;
    assign twf_m0_re[488] = -122;    assign twf_m0_im[488] = 37;
    assign twf_m0_re[489] = -119;    assign twf_m0_im[489] = 48;
    assign twf_m0_re[490] = -114;    assign twf_m0_im[490] = 58;
    assign twf_m0_re[491] = -109;    assign twf_m0_im[491] = 67;
    assign twf_m0_re[492] = -103;    assign twf_m0_im[492] = 76;
    assign twf_m0_re[493] = -96;    assign twf_m0_im[493] = 85;
    assign twf_m0_re[494] = -88;    assign twf_m0_im[494] = 93;
    assign twf_m0_re[495] = -80;    assign twf_m0_im[495] = 100;
    assign twf_m0_re[496] = -71;    assign twf_m0_im[496] = 106;
    assign twf_m0_re[497] = -62;    assign twf_m0_im[497] = 112;
    assign twf_m0_re[498] = -52;    assign twf_m0_im[498] = 117;
    assign twf_m0_re[499] = -42;    assign twf_m0_im[499] = 121;
    assign twf_m0_re[500] = -31;    assign twf_m0_im[500] = 124;
    assign twf_m0_re[501] = -20;    assign twf_m0_im[501] = 126;
    assign twf_m0_re[502] = -9;    assign twf_m0_im[502] = 128;
    assign twf_m0_re[503] = 2;    assign twf_m0_im[503] = 128;
    assign twf_m0_re[504] = 13;    assign twf_m0_im[504] = 127;
    assign twf_m0_re[505] = 23;    assign twf_m0_im[505] = 126;
    assign twf_m0_re[506] = 34;    assign twf_m0_im[506] = 123;
    assign twf_m0_re[507] = 45;    assign twf_m0_im[507] = 120;
    assign twf_m0_re[508] = 55;    assign twf_m0_im[508] = 116;
    assign twf_m0_re[509] = 64;    assign twf_m0_im[509] = 111;
    assign twf_m0_re[510] = 74;    assign twf_m0_im[510] = 105;
    assign twf_m0_re[511] = 82;    assign twf_m0_im[511] = 98;

endmodule
