`timescale 1ns/1ps

module cbfp_mag_detect #(
  parameter DATA_WIDTH = 23, // 입력 비트폭 23비트
  parameter MAG_WIDTH  = $clog2(DATA_WIDTH) + 1 // clog2(23) + 1 = 5 ~ 6 bit : 위치 index 반환용
)(
  input  logic signed [DATA_WIDTH-1:0] din   [15:0], // 16개씩 처리
  output logic        [MAG_WIDTH-1:0]  mag_out [15:0] // 각 입력에 대한 magnitude index 출력
);

  // Case-style leading one detector
  function automatic [MAG_WIDTH-1:0] leading_one(input logic signed [DATA_WIDTH-1:0] val); // 함수: MSB 1의 위치 찾기
    logic [DATA_WIDTH-1:0] abs_val;
    abs_val = val[DATA_WIDTH-1] ? -val : val; 
    // 23비트 입력을 절대값으로 변환 : signed 숫자의 MSB가 1(부호비트 1)이면 음수이므로 부호변환

    // critical path 우려되므로 casez 사용
    casez (abs_val)
      23'b1??????????????????????: return 22;  // MSB가 1인 위치가 22번째, 나머지 don't care
      23'b01?????????????????????: return 21;
      23'b001????????????????????: return 20;
      23'b0001???????????????????: return 19;
      23'b00001??????????????????: return 18;
      23'b000001?????????????????: return 17;
      23'b0000001????????????????: return 16;
      23'b00000001???????????????: return 15;
      23'b000000001??????????????: return 14;
      23'b0000000001?????????????: return 13;
      23'b00000000001????????????: return 12;
      23'b000000000001???????????: return 11;
      23'b0000000000001??????????: return 10;
      23'b00000000000001?????????: return 9;
      23'b000000000000001????????: return 8;
      23'b0000000000000001???????: return 7;
      23'b00000000000000001??????: return 6;
      23'b000000000000000001?????: return 5;
      23'b0000000000000000001????: return 4;
      23'b00000000000000000001???: return 3;
      23'b000000000000000000001??: return 2;
      23'b0000000000000000000001?: return 1;
      23'b00000000000000000000001: return 0;
      default: return 0;
    endcase
  endfunction

  // 16개의 입력에 대해 병렬 처리
  genvar i;
  generate // 하드웨어 반복 구조 자동 생성
    for (i = 0; i < 16; i++) begin : MAG_DET // 1clk 16개 입력에 대해 클럭당 16개씩 detect 처리
      always_comb begin
        mag_out[i] = leading_one(din[i]);
      end
    end
  endgenerate

endmodule
